LIBRARY IEEE;

USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY medicine IS 
	PORT(PULSE: IN STD_LOGIC; 
		CLR: IN STD_LOGIC;
		QD: IN STD_LOGIC; 
		CHECK: IN STD_LOGIC;
		CLK: IN STD_LOGIC;
		CP2: IN STD_LOGIC;
		CP3: IN STD_LOGIC;
		K: IN STD_LOGIC_VECTOR(7 DOWNTO 0);
		DIGIT2,DIGIT3,DIGIT4,DIGIT5: OUT STD_LOGIC_VECTOR(3 DOWNTO 0);
		RED,YELLOW,GREEN: OUT STD_LOGIC;
		MUSIC:OUT STD_LOGIC);
END ENTITY;
	
ARCHITECTURE main OF medicine IS
	
	COMPONENT countclip IS
	PORT(CLIPMAX: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		 CP,CLR: IN STD_LOGIC;
		 CLIPNUMS:OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		 BOTTLENUMS:OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		 TOTAL: OUT STD_LOGIC_VECTOR (11 DOWNTO 0));
	END COMPONENT;
	
	COMPONENT TONES8 IS
	PORT(CP:IN STD_LOGIC;
		 KIND: IN STD_LOGIC;
		 Z:OUT STD_LOGIC);
	END COMPONENT;
	
	SIGNAL EN_FEN,CLR_CLIP,TONES: STD_LOGIC;
	SIGNAL STATE: STD_LOGIC_VECTOR(2 DOWNTO 0):="000";
	SIGNAL BOTTLE, SET_BOTTLE, CURRENT_BOTTLE, FLASH: STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
	SIGNAL CLIP, SET_CLIP, CURRENT_CLIP: STD_LOGIC_VECTOR(7 DOWNTO 0):="00000000";
	SIGNAL TOTAL_CLIP:STD_LOGIC_VECTOR(11 DOWNTO 0):="000000000000";
	
	BEGIN	
		FLASH <= "11111111" WHEN CP3 = '1' ELSE "00000000";
		PROCESS(CLK, FLASH, CP3)
		BEGIN
		IF  RISING_EDGE(CLK) THEN
			CASE STATE IS 
			WHEN "000" => 	
				EN_FEN <= '0';
				SET_BOTTLE <= "00000000";
				SET_CLIP <= "00000000";
				BOTTLE <= "00000000";
				CLIP <= "00000000";
				RED <= '1';
				YELLOW <= '0';
				GREEN <= '0';
				TONES<='0';
			WHEN "001" => 
				EN_FEN <= '0';
				SET_CLIP <= K;
				CLIP <= (K OR FLASH);
				RED <= '0';
				YELLOW <= CP3;
				GREEN <= '0';
			WHEN "010" =>
				EN_FEN <= '1';
				CLR_CLIP<='1';
				SET_BOTTLE <= K;
				CLIP <= SET_CLIP;
				BOTTLE <= (K OR FLASH);
				RED <= '0';
				YELLOW <= CP3;
				GREEN <= '0';
			WHEN "100" =>
				IF CURRENT_BOTTLE = SET_BOTTLE THEN
					EN_FEN <= '0';
					CLR_CLIP<='0';
					CLIP <= SET_CLIP;
					BOTTLE <= SET_BOTTLE;
					RED <= '0';
					YELLOW <= '0';
					GREEN <= '1';
					TONES<='1';
				ELSIF PULSE = '0' THEN
					EN_FEN <= '1';
					CLR_CLIP<='0';
					CLIP <= CURRENT_CLIP;
					BOTTLE <= CURRENT_BOTTLE;
					RED <= '0';
					YELLOW <= '0';
					GREEN <= CP3;
				ELSE
					EN_FEN <= '0';
					CLR_CLIP<='0';
					CLIP <= CURRENT_CLIP;
					BOTTLE <= CURRENT_BOTTLE;
					RED <= '1';
					YELLOW <= '0';
					GREEN <= CP3;
				END IF;
			WHEN "110" =>
				IF CURRENT_BOTTLE = SET_BOTTLE THEN
					EN_FEN <= '0';
					CLR_CLIP <= '0';
					CLIP <= SET_CLIP;
					BOTTLE <= SET_BOTTLE;
					RED <= '0';
					YELLOW <= '0';
					GREEN <= '1';
					TONES<='1';
				ELSIF PULSE = '0' THEN
					EN_FEN <= '1';
					CLR_CLIP<='0';
					CLIP <= SET_CLIP;
					BOTTLE <= SET_BOTTLE;
					RED <= '0';
					YELLOW <= CP3;
					GREEN <= CP3;
				ELSE
					EN_FEN <= '0';
					CLR_CLIP<='0';
					CLIP <= SET_CLIP;
					BOTTLE <= SET_BOTTLE;
					RED <= '1';
					YELLOW <= CP3;
					GREEN <= CP3;
				END IF;			
			WHEN "011" =>
				EN_FEN <= '0';
				CLIP <= (SET_CLIP OR FLASH);
				BOTTLE <= (SET_BOTTLE OR FLASH);
				RED <= CP3;
				YELLOW <= '1';
				GREEN <= '0';
				TONES<='1';
			WHEN OTHERS =>
				
			END CASE;
		END IF;	
		END PROCESS;
	 
		PROCESS (QD, CLR)
		BEGIN
		
		IF CLR = '1' THEN
			STATE <= "000";	
		ELSIF RISING_EDGE(QD) THEN
				CASE STATE IS 
					WHEN "000" => 
						STATE <= "001";
					
					WHEN "001" => 
						STATE <= "010";
					
					WHEN "010" =>
						IF SET_CLIP > "01010000" OR SET_BOTTLE > "00011001" OR SET_CLIP(3 DOWNTO 0) > "1001" OR SET_CLIP(7 DOWNTO 4) > "1001" OR SET_BOTTLE(3 DOWNTO 0) > "1001" OR SET_BOTTLE(7 DOWNTO 4) > "1001" THEN	
							STATE <= "011";
						ELSE
							STATE <= "100";	
						END IF;
						
					WHEN "100" =>
						IF CURRENT_BOTTLE = SET_BOTTLE THEN
							STATE <= "000";
						ELSE
							STATE <= "110";
						END IF;
		
					WHEN "011" =>
						STATE <= "000";
					
					WHEN "110" =>
						IF CURRENT_BOTTLE = SET_BOTTLE THEN
							STATE <= "000";
						ELSE
							STATE <= "100";
						END IF;
				
					WHEN OTHERS =>
						STATE <= "000";
				END CASE;
		END IF;
		
		END PROCESS;
		DIGIT2 <= CLIP(3 DOWNTO 0) WHEN CHECK = '0' ELSE TOTAL_CLIP(3 DOWNTO 0);
		DIGIT3 <= CLIP(7 DOWNTO 4) WHEN CHECK = '0' ELSE TOTAL_CLIP(7 DOWNTO 4);
		DIGIT4 <= BOTTLE(3 DOWNTO 0) WHEN CHECK = '0' ELSE TOTAL_CLIP(11 DOWNTO 8);
		DIGIT5 <= BOTTLE(7 DOWNTO 4) WHEN CHECK = '0' ELSE "ZZZZ";
		cclip: countclip PORT MAP(CLIPMAX=>SET_CLIP,CP=>(CP3 AND EN_FEN),CLR=>CLR_CLIP,CLIPNUMS=>CURRENT_CLIP,BOTTLENUMS=>CURRENT_BOTTLE, TOTAL=>TOTAL_CLIP);
		mu:TONES8 PORT MAP(CP=>(CP2 AND TONES),KIND =>(CP3 AND TONES),Z=>MUSIC);
	END ARCHITECTURE;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY countclip IS
	PORT(CLIPMAX: IN STD_LOGIC_VECTOR (7 DOWNTO 0);
		 CP,CLR: IN STD_LOGIC;
		 CLIPNUMS:OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		 BOTTLENUMS:OUT STD_LOGIC_VECTOR (7 DOWNTO 0);
		 TOTAL: OUT STD_LOGIC_VECTOR (11 DOWNTO 0));
END;
ARCHITECTURE MODE OF countclip IS
	SIGNAL CLIPNUM:STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL BOTTLENUM:STD_LOGIC_VECTOR (7 DOWNTO 0);
	SIGNAL TOTALNUM:STD_LOGIC_VECTOR (11 DOWNTO 0);
	BEGIN
		PROCESS(CP, CLR)
		BEGIN
			IF (CLR = '1') THEN
				CLIPNUM<="00000000";
				BOTTLENUM<="00000000";
				TOTALNUM <="000000000000";
			ELSIF  RISING_EDGE(CP) THEN
				IF TOTALNUM(3 DOWNTO 0)<"1001" THEN 
					TOTALNUM(3 DOWNTO 0)<=TOTALNUM(3 DOWNTO 0)+1;
				ELSE
					TOTALNUM(3 DOWNTO 0)<="0000";
					TOTALNUM(7 DOWNTO 4)<=TOTALNUM(7 DOWNTO 4)+1;
					IF TOTALNUM(7 DOWNTO 4)="1001" THEN
						TOTALNUM(7 DOWNTO 4)<="0000";
						TOTALNUM(11 DOWNTO 8)<=TOTALNUM(11 DOWNTO 8)+1;
					END IF;
						
					IF TOTALNUM(11 DOWNTO 8)="1001" THEN
						TOTALNUM(11 DOWNTO 8)<="0000";
						TOTALNUM(7 DOWNTO 4)<="0000";
						TOTALNUM(3 DOWNTO 0)<="0000";
					END IF;
				END IF;
					
				IF (CLIPNUM=CLIPMAX) THEN
					IF (BOTTLENUM(3 DOWNTO 0)="1001") THEN
						BOTTLENUM(3 DOWNTO 0)<="0000";
						BOTTLENUM(7 DOWNTO 4)<=BOTTLENUM(7 DOWNTO 4) + 1;
					ELSE
						BOTTLENUM(3 DOWNTO 0)<=BOTTLENUM(3 DOWNTO 0) + 1;
					END IF;
					CLIPNUM<="00000001";
				ELSIF (CLIPNUM(3 DOWNTO 0)="1001") THEN
					CLIPNUM(3 DOWNTO 0)<="0000";
					CLIPNUM(7 DOWNTO 4)<=CLIPNUM(7 DOWNTO 4) + 1;
				ELSE
					CLIPNUM(3 DOWNTO 0)<=CLIPNUM(3 DOWNTO 0) + 1;		
				END IF;
			END IF;
		END PROCESS;
		CLIPNUMS<=CLIPNUM;
		BOTTLENUMS<=BOTTLENUM;
		TOTAL<=TOTALNUM;
END MODE;

LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY TONES8 IS
	PORT(CP:IN STD_LOGIC;
		 KIND: IN STD_LOGIC;
		 Z:OUT STD_LOGIC);
END;
ARCHITECTURE SPKOUT OF TONES8 IS
	SIGNAL COUNT:STD_LOGIC_VECTOR(1 DOWNTO 0);
	SIGNAL STA:STD_LOGIC;
	BEGIN	
		PROCESS(CP)
		BEGIN
			IF RISING_EDGE(CP) THEN
				IF (COUNT="11") THEN
					COUNT<="00";
					STA <= NOT STA;
				ELSE
					COUNT<=COUNT+1;
				END IF;
			END IF;
		END PROCESS;
		Z <= CP WHEN KIND = '0' ELSE STA;
END SPKOUT;