LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY control IS
	PORT(CP_QD, CLOCK, ALARM,CP_CM,CP_AH,CP_AM, CP: IN STD_LOGIC;
		SET_OUT: OUT STD_LOGIC;
		SET_M:OUT STD_LOGIC_VECTOR(2 DOWNTO 0));
END ENTITY;

ARCHITECTURE control_func OF control IS
	SIGNAL SET: STD_LOGIC:='0'; 
	SIGNAL SET_MODE: STD_LOGIC_VECTOR(2 DOWNTO 0):="000";
	BEGIN
	
	SET <= '1' WHEN (CLOCK = '1' OR ALARM = '1') ELSE '0';
	
	PROCESS (CP_QD, SET)
	BEGIN
		IF SET = '0' THEN
			SET_MODE <= "000";
		ELSIF RISING_EDGE(CP_QD) THEN 
			IF SET_MODE = "000" THEN
				SET_MODE <= "001";
			END IF;
				
			CASE SET_MODE IS
				WHEN "001" => SET_MODE <= "010";
				WHEN "010" => SET_MODE <= "100";
				WHEN "100" => SET_MODE <= "001";
				WHEN OTHERS => SET_MODE <= "001";
			END CASE;
		END IF;
	END PROCESS;
	
	SET_M <= SET_MODE;
	SET_OUT <= SET;
END ARCHITECTURE;