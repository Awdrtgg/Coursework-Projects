LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.STD_LOGIC_UNSIGNED.ALL;

ENTITY decoder IS
	PORT(INPUT: IN STD_LOGIC_VECTOR(3 DOWNTO 0);
		OUTPUT:OUT STD_LOGIC_VECTOR(6 DOWNTO 0));
END ENTITY;

ARCHITECTURE decoder_func OF decoder IS
	BEGIN
	OUTPUT <= 	"0111111" WHEN INPUT = "0000" ELSE
				"0000110" WHEN INPUT = "0001" ELSE
				"1011011" WHEN INPUT = "0010" ELSE
				"1001111" WHEN INPUT = "0011" ELSE
				"1100110" WHEN INPUT = "0100" ELSE
				"1101101" WHEN INPUT = "0101" ELSE
				"1111101" WHEN INPUT = "0110" ELSE
				"0000111" WHEN INPUT = "0111" ELSE
				"1111111" WHEN INPUT = "1000" ELSE
				"1101111" WHEN INPUT = "1001" ELSE
								"0000000";
END ARCHITECTURE;